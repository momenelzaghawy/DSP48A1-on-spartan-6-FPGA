module DSP48A1 (CLK,OPMODE,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP,RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,BCOUT,PCIN,PCOUT,A,B,C,D,CARRYIN,M,P,CARRYOUT,CARRYOUTF,BCIN);
parameter A0REG=0,A1REG=1,B0REG=0,B1REG=1,CREG=1,DREG=1,MREG=1,PREG=1,CARRYINREG=1,CARRYOUTREG=1,OPMODEREG=1;
parameter CARRYINSEL=1,B_INPUT=1,RSTTYPE="SYNC";
input [17:0]A,B,D,BCIN;
input [47:0]C,PCIN;
input CARRYIN,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP;
input RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,CLK;
input [7:0]OPMODE;
output [35:0]M;
output [47:0]P,PCOUT;
output [17:0]BCOUT;
output CARRYOUT,CARRYOUTF;
wire [17:0]D_w,A_w,B_mux,B_w,add_sub1,add_sub1_w,B1_reg_w,A1_reg_w;
wire [47:0]C_w,mux_x,mux_z,add_sub2_w,P_w;
wire [35:0]mult_w,mult1_w;
wire [7:0]OPMODE_w;
wire carryin0_w,CIN,carry_w,CARRYOUT_reg;
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(DREG),.N(18)) D0 (.d(D),.CLK(CLK),.RST(RSTD),.E(CED),.q(D_w));
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(A0REG),.N(18)) A0 (.d(A),.CLK(CLK),.RST(RSTA),.E(CEA),.q(A_w));
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(CREG),.N(48)) C0 (.d(C),.CLK(CLK),.RST(RSTC),.E(CEC),.q(C_w));
assign B_mux=(B_INPUT==1)? B :(B_INPUT==0)? BCIN : 0;
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(B0REG),.N(18)) B0 (.d(B_mux),.CLK(CLK),.RST(RSTB),.E(CEB),.q(B_w));
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(OPMODEREG),.N(8)) opmode0 (.d(OPMODE),.CLK(CLK),.RST(RSTOPMODE),.E(CEOPMODE),.q(OPMODE_w));
assign add_sub1=(OPMODE_w[6]==0)? (D_w + B_w) : (D_w - B_w);
assign add_sub1_w=(OPMODE_w[4]==0)? B_w : add_sub1;  
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(B1REG),.N(18)) B1 (.d(add_sub1_w),.CLK(CLK),.RST(RSTB),.E(CEB),.q(B1_reg_w));
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(A1REG),.N(18)) A1 (.d(A_w),.CLK(CLK),.RST(RSTA),.E(CEA),.q(A1_reg_w));
assign mult_w=A1_reg_w * B1_reg_w ;
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(MREG),.N(36)) M0 (.d(mult_w),.CLK(CLK),.RST(RSTM),.E(CEM),.q(mult1_w));
assign M=mult1_w;
assign mux_x=(OPMODE_w[1:0]==0)? 0 :(OPMODE_w[1:0]==1)? {12'b0,mult1_w} : (OPMODE_w[1:0]==2)? P_w : {D_w[11:0],A1_reg_w[17:0],B1_reg_w[17:0]};
assign mux_z=(OPMODE_w[3:2]==0)? 0 :(OPMODE_w[3:2]==1)? PCIN : (OPMODE_w[3:2]==2)? P_w : C_w ;
assign carryin0_w=(CARRYINSEL==1)? OPMODE_w[5] : (CARRYINSEL==0)? CARRYIN : 0;
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(CARRYINREG),.N(1)) carryin0 (.d(carryin0_w),.CLK(CLK),.RST(RSTCARRYIN),.E(CECARRYIN),.q(CIN));
assign {carry_w,add_sub2_w}=(OPMODE_w[7]==0)? mux_z+mux_x+CIN : mux_z - (mux_x + CIN);
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(PREG),.N(48)) P0 (.d(add_sub2_w),.CLK(CLK),.RST(RSTP),.E(CEP),.q(P_w));
assign P=P_w;
assign PCOUT=P_w;
reg_mux #(.RSTTYPE(RSTTYPE),.PYPLINE(CARRYOUTREG),.N(1)) cout0 (.d(carry_w),.CLK(CLK),.RST(RSTCARRYIN),.E(CECARRYIN),.q(CARRYOUT_reg));
assign CARRYOUT=CARRYOUT_reg;
assign CARRYOUTF=CARRYOUT_reg;
assign BCOUT=B1_reg_w;
endmodule